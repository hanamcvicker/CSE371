// The inputs are the clock and reset provided by DE1-SoC, and outer and inner, the sensor inputs. 
// The output is count, which holds the number of cars currently in the lot.

module parking_lot_occupancy (clk, reset, count, outer, inner);

	input logic clk, reset, outer, inner;
	logic enter, exit;
	
	output logic [4:0] count;
	
	logic outerq;
	double_FF outerFF (.q(outerq), .d(outer), .reset, .clk);
	logic innerq;
	double_FF innerFF (.q(innerq), .d(inner), .reset, .clk);
	
	carDetect cd (.clk, .reset, .outer(outerq), .inner(innerq), .enter, .exit);
	car_counter cc (.clk, .reset, .incr(enter), .decr(exit), .count);
	

endmodule

module parking_lot_occupancy_testbench();  
	logic  clk, reset, outer, inner;  
	logic  [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;  
  
	parking_lot_occupancy dut (clk, reset, outer, inner, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5);   
   
	// Set up a simulated clock.   
	parameter CLOCK_PERIOD=100;  
	initial begin  
		clk <= 0;  
		forever #(CLOCK_PERIOD/2) clk <= ~clk; // Forever toggle the clock 
	end  
   
 initial begin  
															@(posedge clk);   
  reset <= 1;         								@(posedge clk);  
  reset <= 0; outer <= 0; inner <= 0; 			@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
  outer <= 1; 											@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
  inner <= 1; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
  outer <= 0; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
  inner <= 0; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
  outer <= 1; 									   	@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
  inner <= 1; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
  outer <= 0; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
  inner <= 0; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
  outer <= 1; 											@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
  inner <= 1; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   inner <= 1; 										@(posedge clk);   
													      @(posedge clk);   
														   @(posedge clk);   
    outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	 inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
    outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
    inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
    outer <= 0;										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	 inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
    outer <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
    inner <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
    outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	 inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	 inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
    outer <= 1;										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
    inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	 outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
   inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
	inner <= 1;											@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
	inner <= 1;											@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   inner <= 1;											@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0;											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
   inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);  
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
	inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
  inner <= 0; 											@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
	outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk); 
   inner <= 1; 										@(posedge clk);
															@(posedge clk);
															@(posedge clk);			 
   outer <= 1; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);   
   inner <= 0; 										@(posedge clk);   
															@(posedge clk);   
															@(posedge clk);
   outer <= 0; 										@(posedge clk);   
															@(posedge clk);   
                    
	
  $stop; // End the simulation.  
 end  
endmodule  